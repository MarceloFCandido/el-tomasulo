module instrQueue();
	
endmodule
