module multiplexador(Entrada1, Entrada2, Entrada3, Entrada4, Seletor, Saida); 



endmodule
