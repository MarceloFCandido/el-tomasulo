module CDB_Arbt(UA_as, UA_ls, Un_mem, CDB);	//Recebe as saidas das UF's e decide qual ira para o CDB
	



endmodule
